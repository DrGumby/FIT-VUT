library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;
use std.textio.all;

-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity testbench is
end entity testbench;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture behavioral of testbench is

   signal smclk   : std_logic := '1';
   signal aclk    : std_logic;
   signal fclk    : std_logic;

   signal ledf  : std_logic;
   signal p3m   : std_logic_vector(7 downto 0) := (others=>'Z');   
   signal afbus : std_logic_vector(11 downto 0) :=(others =>'Z');
   signal xbus  : std_logic_vector(45 downto 0) :=(others =>'Z');
   signal rdbus : std_logic_vector(7 downto 0) :=(others =>'Z');
   signal ldbus : std_logic_vector(7 downto 0) :=(others =>'Z');

   signal ispi_clk : std_logic:='1';
   signal ispi_cs  : std_logic:='1';
   signal ispi_di  : std_logic:='Z';    
   signal ispi_do  : std_logic:='1';
   
begin
   --Unit under test
   uut: entity work.fpga
      port map(
         SMCLK    => smclk,
         ACLK    => aclk,
         FCLK    => fclk,
         LEDF     => ledf,
   
         SPI_CLK  => ispi_clk,
         SPI_CS   => '1',
         SPI_FPGA_CS => ispi_cs,
         SPI_DI   => ispi_di,
         SPI_DO   => ispi_do,
   
         KIN      => open,
         KOUT     => (others => 'Z'),
   
         LE       => open,
         LRW      => open,
         LRS      => open,
         LD       => ldbus,

         RA       => open,
         RD       => rdbus,
         RDQM     => open,
         RCS      => open,
         RRAS     => open,
         RCAS     => open,
         RWE      => open,
         RCKE     => open,
         RCLK     => open,

         P3M      => p3m,
         AFBUS    => afbus,
   	   X        => xbus
   );

   -- Clock generator (SMCLK) 7.3725 MHz
   smclk <= not smclk after 67.819 ns;
	
   
   -- SPI clock generator (SMCLK/4)
   ispi_clk <= not ispi_clk after 271.276 ns;
   
   -- Reset generator
   p3m(0) <= '1', '0' after 1000 ns;

   -- Test bench circuit
   write:process
   begin
      ispi_cs <= '1';
      ispi_di <= 'Z';
      ispi_do <= '1';
      wait until p3m(0)='0';
      wait for 100 ns;

      -- test bench
      wait;
   end process;

end architecture behavioral;

